

constant integer STATE_NONE = 0;
constant integer STATE_RESET = 1;
constant integer STATE_FETCH = 2;
constant integer STATE_DECODE = 3;
constant integer STATE_STORE = 4;


constant integer STATE_HALT = 0xFF;


constant integer VBIT = 3;
constant integer NBIT = 2;
constant integer CBIT = 1;
constant integer ZBIT = 0;

typedef struct
{
   bit[16] value;
} reg_type;

module lsa_core
(
    clock          in_clock,
    input  bit     in_reset
)
{
    default clock in_clock ;
    default reset active_low in_reset ;

    clocked reg_type[64] reg = {{value=0}};

    comb bit[16] pc_next;

    clocked bit[4] astate = STATE_NONE;
    comb bit[4] astate_next;

    clocked bit[16] inst = 0;

    comb bit[17] op_a;
    comb bit[17] op_b;
    comb bit[17] op_res;


    comb bit[16] mem_add;
    comb bit[16] mem_out;
    comb bit[16] mem_in;
    comb bit[1]  mem_wr;
    comb bit[1]  mem_rd;
    comb bit[1]  mem_fetch;

    clocked bit[8] leds = 0x00;


    the_mem:
    {
        mem_out = 0x0000;
        if(mem_rd == 1b1)
        {
            full_switch(mem_add)
            {

case 16h0000: { mem_out = 0xC001; }
case 16h0001: { mem_out = 0xC000; }
case 16h0002: { mem_out = 0x97F1; }
case 16h0003: { mem_out = 0x8500; }
case 16h0004: { mem_out = 0x8820; }
case 16h0005: { mem_out = 0x6889; }
case 16h0006: { mem_out = 0xC2FE; }
case 16h0007: { mem_out = 0x6558; }
case 16h0008: { mem_out = 0x4758; }
case 16h0009: { mem_out = 0x8820; }
case 16h000A: { mem_out = 0xC0FA; }


                default:
                {
                    mem_out = 0x0000;
                }
            }
        }
        if(mem_wr == 1)
        {
            full_switch(mem_add)
            {
                case 0xF100:
                {
                    leds <= mem_in[8;0];
                }
                default:
                {
                }
            }
        }




    }

    the_code:
    {
        mem_add   = 0x0000;
        mem_in    = 0x0000;
        mem_wr    = 0;
        mem_rd    = 0;
        mem_fetch = 0;
        astate_next = astate;
        pc_next = reg[0].value;


        full_switch(astate)
        {
            case STATE_NONE:
            {
                astate_next = STATE_RESET;
            }
            case STATE_RESET:
            {
                pc_next = 0x0000;
                astate_next = STATE_FETCH;
            }
            case STATE_FETCH:
            {
                pc_next = reg[0].value + 1;
                mem_add = reg[0].value;
                mem_fetch = 1;
                mem_rd = 1;
                inst <= mem_out;
                astate_next = STATE_DECODE;
            }
            case STATE_DECODE:
            {
                astate_next = STATE_HALT;
                full_switch(inst[4;12])
                {
                    case 0x4: //0100 dddd ssss aaaa  load/store
                    {
                        full_switch(inst[4;0])
                        {
                            case 0x8: //1000 stw [rd]  ,rs
                            {
                                //1000 stw [rd]  ,rs
                                mem_add = reg[bundle(2b0,inst[4;8])].value;
                                mem_wr = 1;
                                mem_in = reg[bundle(2b0,inst[4;4])].value;
                                astate_next = STATE_STORE;
                            }
                            default:
                            {
                                astate_next = STATE_HALT;
                            }
                        }
                    }
                    case 0x6:
                    {
                        full_switch(inst[4;0])
                        {
                            case 0x8:
                            {
                                //1000 inc rd,rs
                                op_a = 17b1;
                                op_b = bundle(1b0,reg[bundle(2b0,inst[4;4])].value);
                                op_res = op_a + op_b;
                                reg[1].value[CBIT] <= op_res[16];
                                reg[1].value[NBIT] <= op_res[15];

                                if(op_res[16;0] == 16h0000)
                                {
                                    reg[1].value[ZBIT] <= 1b1;
                                }
                                else
                                {
                                    reg[1].value[ZBIT] <= 1b0;
                                }
                                if((op_a[15] == op_b[15]) && (op_res[15] != op_b[15] ) )
                                {
                                    reg[1].value[VBIT] <= 1b1;
                                }
                                else
                                {
                                    reg[1].value[VBIT] <= 1b0;
                                }
                                reg[bundle(2b0,inst[4;8])].value <= op_res[16;0];
                                astate_next = STATE_FETCH;
                            }
                            case 0x9: //dec rd,rd
                            {
                                //1001 dec rd,rs
                                op_a = bundle(1b0,reg[bundle(2b0,inst[4;4])].value);
                                op_b = 17b1;
                                op_res = op_a - op_b;
                                reg[1].value[CBIT] <= (~op_res[16]);
                                reg[1].value[NBIT] <= op_res[15];

                                if(op_res[16;0] == 16h0000)
                                {
                                    reg[1].value[ZBIT] <= 1b1;
                                }
                                else
                                {
                                    reg[1].value[ZBIT] <= 1b0;
                                }
                                if((op_a[15] != op_b[15]) && (op_res[15] == op_b[15] ) )
                                {
                                    reg[1].value[VBIT] <= 1b1;
                                }
                                else
                                {
                                    reg[1].value[VBIT] <= 1b0;
                                }
                                reg[bundle(2b0,inst[4;8])].value <= op_res[16;0];
                                astate_next = STATE_FETCH;

                            }
                            default:
                            {
                                astate_next = STATE_HALT;
                            }
                        }
                    }
                    case 0x8: //llz rd,#imm
                    {
                        reg[bundle(2b00,inst[4;8])].value[8;8] <= 0x00;
                        reg[bundle(2b00,inst[4;8])].value[8;0] <= inst[8;0];
                        astate_next = STATE_FETCH;
                    }
                    case 0x9: //lhz rd,#imm
                    {
                        reg[bundle(2b00,inst[4;8])].value[8;8] <= inst[8;0];
                        reg[bundle(2b00,inst[4;8])].value[8;0] <= 0x00;
                        astate_next = STATE_FETCH;
                    }
                    case 0xA: //ll rd,#imm
                    {
                        reg[bundle(2b00,inst[4;8])].value[8;0] <= inst[8;0];
                        astate_next = STATE_FETCH;
                    }
                    case 0xB: //lh rd,#imm
                    {
                        reg[bundle(2b00,inst[4;8])].value[8;8] <= inst[8;0];
                        astate_next = STATE_FETCH;
                    }
                    case 0xC:
                    {
                        full_switch(inst[4;8])
                        {
                            case 0x0: //b unconditional
                            {
                                pc_next = reg[0].value + bundle(inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[8;0]);
                                astate_next = STATE_FETCH;
                            }
                            case 0x1: //bz
                            {
                                if(reg[1].value[ZBIT] == 1)
                                {
                                    pc_next = reg[0].value + bundle(inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[8;0]);
                                }
                                astate_next = STATE_FETCH;
                            }
                            case 0x2: //bnz
                            {
                                if(reg[1].value[ZBIT] == 0)
                                {
                                    pc_next = reg[0].value + bundle(inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[7],inst[8;0]);
                                }
                                astate_next = STATE_FETCH;
                            }
                            default:
                            {
                                astate_next = STATE_HALT;
                            }
                        }
                    }
                    default:
                    {
                        astate_next = STATE_HALT;
                    }
                }


            }

            case STATE_STORE:
            {
                astate_next = STATE_FETCH;
            }
            default:
            {
                astate_next = STATE_HALT;
            }
        }


        reg[0].value <= pc_next;

        astate <= astate_next;
    }
}
